library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity skutusu is port 
(
	byte : in std_logic_vector(7 downto 0);
	bytecikis : out std_logic_vector(7 downto 0)
);
end skutusu;

architecture degisim of skutusu is

	begin
	process(byte)	
	begin
		case byte is
				when x"00" => bytecikis <= x"63";
				when x"01" => bytecikis <= x"7c";
				when x"02" => bytecikis <= x"77";
				when x"03" => bytecikis <= x"7b";
				when x"04" => bytecikis <= x"f2";
				when x"05" => bytecikis <= x"6b";
				when x"06" => bytecikis <= x"6f";
				when x"07" => bytecikis <= x"c5";
				when x"08" => bytecikis <= x"30";
				when x"09" => bytecikis <= x"01";
				when x"0a" => bytecikis <= x"67";
				when x"0b" => bytecikis <= x"2b";
				when x"0c" => bytecikis <= x"fe";
				when x"0d" => bytecikis <= x"d7";
				when x"0e" => bytecikis <= x"ab";
				when x"0f" => bytecikis <= x"76";
				when x"10" => bytecikis <= x"ca";
				when x"11" => bytecikis <= x"82";
				when x"12" => bytecikis <= x"c9";
				when x"13" => bytecikis <= x"7d";
				when x"14" => bytecikis <= x"fa";
				when x"15" => bytecikis <= x"59";
				when x"16" => bytecikis <= x"47";
				when x"17" => bytecikis <= x"f0";
				when x"18" => bytecikis <= x"ad";
				when x"19" => bytecikis <= x"d4";
				when x"1a" => bytecikis <= x"a2";
				when x"1b" => bytecikis <= x"af";
				when x"1c" => bytecikis <= x"9c";
				when x"1d" => bytecikis <= x"a4";
				when x"1e" => bytecikis <= x"72";
				when x"1f" => bytecikis <= x"c0";
				when x"20" => bytecikis <= x"b7";
				when x"21" => bytecikis <= x"fd";
				when x"22" => bytecikis <= x"93";
				when x"23" => bytecikis <= x"26";
				when x"24" => bytecikis <= x"36";
				when x"25" => bytecikis <= x"3f";
				when x"26" => bytecikis <= x"f7";
				when x"27" => bytecikis <= x"cc";
				when x"28" => bytecikis <= x"34";
				when x"29" => bytecikis <= x"a5";
				when x"2a" => bytecikis <= x"e5";
				when x"2b" => bytecikis <= x"f1";
				when x"2c" => bytecikis <= x"71";
				when x"2d" => bytecikis <= x"d8";
				when x"2e" => bytecikis <= x"31";
				when x"2f" => bytecikis <= x"15";
				when x"30" => bytecikis <= x"04";
				when x"31" => bytecikis <= x"c7";
				when x"32" => bytecikis <= x"23";
				when x"33" => bytecikis <= x"c3";
				when x"34" => bytecikis <= x"18";
				when x"35" => bytecikis <= x"96";
				when x"36" => bytecikis <= x"05";
				when x"37" => bytecikis <= x"9a";
				when x"38" => bytecikis <= x"07";
				when x"39" => bytecikis <= x"12";
				when x"3a" => bytecikis <= x"80";
				when x"3b" => bytecikis <= x"e2";
				when x"3c" => bytecikis <= x"eb";
				when x"3d" => bytecikis <= x"27";
				when x"3e" => bytecikis <= x"b2";
				when x"3f" => bytecikis <= x"75";
				when x"40" => bytecikis <= x"09";
				when x"41" => bytecikis <= x"83";
				when x"42" => bytecikis <= x"2c";
				when x"43" => bytecikis <= x"1a";
				when x"44" => bytecikis <= x"1b";
				when x"45" => bytecikis <= x"6e";
				when x"46" => bytecikis <= x"5a";
				when x"47" => bytecikis <= x"a0";
				when x"48" => bytecikis <= x"52";
				when x"49" => bytecikis <= x"3b";
				when x"4a" => bytecikis <= x"d6";
				when x"4b" => bytecikis <= x"b3";
				when x"4c" => bytecikis <= x"29";
				when x"4d" => bytecikis <= x"e3";
				when x"4e" => bytecikis <= x"2f";
				when x"4f" => bytecikis <= x"84";
				when x"50" => bytecikis <= x"53";
				when x"51" => bytecikis <= x"d1";
				when x"52" => bytecikis <= x"00";
				when x"53" => bytecikis <= x"ed";
				when x"54" => bytecikis <= x"20";
				when x"55" => bytecikis <= x"fc";
				when x"56" => bytecikis <= x"b1";
				when x"57" => bytecikis <= x"5b";
				when x"58" => bytecikis <= x"6a";
				when x"59" => bytecikis <= x"cb";
				when x"5a" => bytecikis <= x"be";
				when x"5b" => bytecikis <= x"39";
				when x"5c" => bytecikis <= x"4a";
				when x"5d" => bytecikis <= x"4c";
				when x"5e" => bytecikis <= x"58";
				when x"5f" => bytecikis <= x"cf";
				when x"60" => bytecikis <= x"d0";
				when x"61" => bytecikis <= x"ef";
				when x"62" => bytecikis <= x"aa";
				when x"63" => bytecikis <= x"fb";
				when x"64" => bytecikis <= x"43";
				when x"65" => bytecikis <= x"4d";
				when x"66" => bytecikis <= x"33";
				when x"67" => bytecikis <= x"85";
				when x"68" => bytecikis <= x"45";
				when x"69" => bytecikis <= x"f9";
				when x"6a" => bytecikis <= x"02";
				when x"6b" => bytecikis <= x"7f";
				when x"6c" => bytecikis <= x"50";
				when x"6d" => bytecikis <= x"3c";
				when x"6e" => bytecikis <= x"9f";
				when x"6f" => bytecikis <= x"a8";
				when x"70" => bytecikis <= x"51";
				when x"71" => bytecikis <= x"a3";
				when x"72" => bytecikis <= x"40";
				when x"73" => bytecikis <= x"8f";
				when x"74" => bytecikis <= x"92";
				when x"75" => bytecikis <= x"9d";
				when x"76" => bytecikis <= x"38";
				when x"77" => bytecikis <= x"f5";
				when x"78" => bytecikis <= x"bc";
				when x"79" => bytecikis <= x"b6";
				when x"7a" => bytecikis <= x"da";
				when x"7b" => bytecikis <= x"21";
				when x"7c" => bytecikis <= x"10";
				when x"7d" => bytecikis <= x"ff";
				when x"7e" => bytecikis <= x"f3";
				when x"7f" => bytecikis <= x"d2";
				when x"80" => bytecikis <= x"cd";
				when x"81" => bytecikis <= x"0c";
				when x"82" => bytecikis <= x"13";
				when x"83" => bytecikis <= x"ec";
				when x"84" => bytecikis <= x"5f";
				when x"85" => bytecikis <= x"97";
				when x"86" => bytecikis <= x"44";
				when x"87" => bytecikis <= x"17";
				when x"88" => bytecikis <= x"c4";
				when x"89" => bytecikis <= x"a7";
				when x"8a" => bytecikis <= x"7e";
				when x"8b" => bytecikis <= x"3d";
				when x"8c" => bytecikis <= x"64";
				when x"8d" => bytecikis <= x"5d";
				when x"8e" => bytecikis <= x"19";
				when x"8f" => bytecikis <= x"73";
				when x"90" => bytecikis <= x"60";
				when x"91" => bytecikis <= x"81";
				when x"92" => bytecikis <= x"4f";
				when x"93" => bytecikis <= x"dc";
				when x"94" => bytecikis <= x"22";
				when x"95" => bytecikis <= x"2a";
				when x"96" => bytecikis <= x"90";
				when x"97" => bytecikis <= x"88";
				when x"98" => bytecikis <= x"46";
				when x"99" => bytecikis <= x"ee";
				when x"9a" => bytecikis <= x"b8";
				when x"9b" => bytecikis <= x"14";
				when x"9c" => bytecikis <= x"de";
				when x"9d" => bytecikis <= x"5e";
				when x"9e" => bytecikis <= x"0b";
				when x"9f" => bytecikis <= x"db";
				when x"a0" => bytecikis <= x"e0";
				when x"a1" => bytecikis <= x"32";
				when x"a2" => bytecikis <= x"3a";
				when x"a3" => bytecikis <= x"0a";
				when x"a4" => bytecikis <= x"49";
				when x"a5" => bytecikis <= x"06";
				when x"a6" => bytecikis <= x"24";
				when x"a7" => bytecikis <= x"5c";
				when x"a8" => bytecikis <= x"c2";
				when x"a9" => bytecikis <= x"d3";
				when x"aa" => bytecikis <= x"ac";
				when x"ab" => bytecikis <= x"62";
				when x"ac" => bytecikis <= x"91";
				when x"ad" => bytecikis <= x"95";
				when x"ae" => bytecikis <= x"e4";
				when x"af" => bytecikis <= x"79";
				when x"b0" => bytecikis <= x"e7";
				when x"b1" => bytecikis <= x"c8";
				when x"b2" => bytecikis <= x"37";
				when x"b3" => bytecikis <= x"6d";
				when x"b4" => bytecikis <= x"8d";
				when x"b5" => bytecikis <= x"d5";
				when x"b6" => bytecikis <= x"4e";
				when x"b7" => bytecikis <= x"a9";
				when x"b8" => bytecikis <= x"6c";
				when x"b9" => bytecikis <= x"56";
				when x"ba" => bytecikis <= x"f4";
				when x"bb" => bytecikis <= x"ea";
				when x"bc" => bytecikis <= x"65";
				when x"bd" => bytecikis <= x"7a";
				when x"be" => bytecikis <= x"ae";
				when x"bf" => bytecikis <= x"08";
				when x"c0" => bytecikis <= x"ba";
				when x"c1" => bytecikis <= x"78";
				when x"c2" => bytecikis <= x"25";
				when x"c3" => bytecikis <= x"2e";
				when x"c4" => bytecikis <= x"1c";
				when x"c5" => bytecikis <= x"a6";
				when x"c6" => bytecikis <= x"b4";
				when x"c7" => bytecikis <= x"c6";
				when x"c8" => bytecikis <= x"e8";
				when x"c9" => bytecikis <= x"dd";
				when x"ca" => bytecikis <= x"74";
				when x"cb" => bytecikis <= x"1f";
				when x"cc" => bytecikis <= x"4b";
				when x"cd" => bytecikis <= x"bd";
				when x"ce" => bytecikis <= x"8b";
				when x"cf" => bytecikis <= x"8a";
				when x"d0" => bytecikis <= x"70";
				when x"d1" => bytecikis <= x"3e";
				when x"d2" => bytecikis <= x"b5";
				when x"d3" => bytecikis <= x"66";
				when x"d4" => bytecikis <= x"48";
				when x"d5" => bytecikis <= x"03";
				when x"d6" => bytecikis <= x"f6";
				when x"d7" => bytecikis <= x"0e";
				when x"d8" => bytecikis <= x"61";
				when x"d9" => bytecikis <= x"35";
				when x"da" => bytecikis <= x"57";
				when x"db" => bytecikis <= x"b9";
				when x"dc" => bytecikis <= x"86";
				when x"dd" => bytecikis <= x"c1";
				when x"de" => bytecikis <= x"1d";
				when x"df" => bytecikis <= x"9e";
				when x"e0" => bytecikis <= x"e1";
				when x"e1" => bytecikis <= x"f8";
				when x"e2" => bytecikis <= x"98";
				when x"e3" => bytecikis <= x"11";
				when x"e4" => bytecikis <= x"69";
				when x"e5" => bytecikis <= x"d9";
				when x"e6" => bytecikis <= x"8e";
				when x"e7" => bytecikis <= x"94";
				when x"e8" => bytecikis <= x"9b";
				when x"e9" => bytecikis <= x"1e";
				when x"ea" => bytecikis <= x"87";
				when x"eb" => bytecikis <= x"e9";
				when x"ec" => bytecikis <= x"ce";
				when x"ed" => bytecikis <= x"55";
				when x"ee" => bytecikis <= x"28";
				when x"ef" => bytecikis <= x"df";
				when x"f0" => bytecikis <= x"8c";
				when x"f1" => bytecikis <= x"a1";
				when x"f2" => bytecikis <= x"89";
				when x"f3" => bytecikis <= x"0d";
				when x"f4" => bytecikis <= x"bf";
				when x"f5" => bytecikis <= x"e6";
				when x"f6" => bytecikis <= x"42";
				when x"f7" => bytecikis <= x"68";
				when x"f8" => bytecikis <= x"41";
				when x"f9" => bytecikis <= x"99";
				when x"fa" => bytecikis <= x"2d";
				when x"fb" => bytecikis <= x"0f";
				when x"fc" => bytecikis <= x"b0";
				when x"fd" => bytecikis <= x"54";
				when x"fe" => bytecikis <= x"bb";
				when x"ff" => bytecikis <= x"16";			
				when others=> bytecikis <= x"00";
		end case;
	end process;
end degisim;